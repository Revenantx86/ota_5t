* Extracted by KLayout with SKY130 LVS runset on : 29/08/2024 17:10

.SUBCKT ota_5t
M$1 \$7 \$7 VDD \$9 sky130_fd_pr__pfet_01v8 L=1 W=1.5 AS=0.45 AD=0.375 PS=3.6
+ PD=2
M$2 VDD \$7 \$7 \$9 sky130_fd_pr__pfet_01v8 L=1 W=1.5 AS=0.375 AD=0.375 PS=2
+ PD=2
M$3 \$7 \$7 VDD \$9 sky130_fd_pr__pfet_01v8 L=1 W=1.5 AS=0.375 AD=0.45 PS=2
+ PD=3.6
M$4 Vout \$7 VDD \$9 sky130_fd_pr__pfet_01v8 L=1 W=1.5 AS=0.45 AD=0.375 PS=3.6
+ PD=2
M$5 VDD \$7 Vout \$9 sky130_fd_pr__pfet_01v8 L=1 W=1.5 AS=0.375 AD=0.375 PS=2
+ PD=2
M$6 Vout \$7 VDD \$9 sky130_fd_pr__pfet_01v8 L=1 W=1.5 AS=0.375 AD=0.45 PS=2
+ PD=3.6
M$7 \$5 Vn Vout sky130_gnd sky130_fd_pr__nfet_01v8 L=0.5 W=3 AS=0.9 AD=0.9
+ PS=6.6 PD=6.6
M$8 \$5 Vp \$7 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.5 W=3 AS=0.9 AD=0.9
+ PS=6.6 PD=6.6
M$9 VSS Ib \$5 sky130_gnd sky130_fd_pr__nfet_01v8 L=1 W=4 AS=1.2 AD=1.2 PS=8.6
+ PD=8.6
M$10 Ib Ib VSS sky130_gnd sky130_fd_pr__nfet_01v8 L=1 W=4 AS=1.2 AD=1.2 PS=8.6
+ PD=8.6
.ENDS ota_5t
