* NGSPICE file created from ota_5t.ext - technology: sky130A

.subckt ota_5t Ib Vn Vp Vout VDD VSS
X0 VDD.t7 a_2521_2520.t3 a_2521_2520.t4 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.375 pd=2 as=0.45 ps=3.6 w=1.5 l=1
X1 a_2521_2520.t0 Vp.t0 a_2521_2360# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.9 pd=6.6 as=0.9 ps=6.6 w=3 l=0.5
X2 a_2521_2520.t6 a_2521_2520.t5 VDD.t6 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.375 pd=2 as=0.375 ps=2 w=1.5 l=1
X3 Vout.t0 Vn.t0 a_2521_2360# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.9 pd=6.6 as=0.9 ps=6.6 w=3 l=0.5
X4 VDD.t5 a_2521_2520.t1 a_2521_2520.t2 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.6 as=0.375 ps=2 w=1.5 l=1
X5 VSS.t1 Ib.t0 Ib.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=1.2 ps=8.6 w=4 l=1
X6 VDD.t3 a_2521_2520.t7 Vout.t3 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.375 pd=2 as=0.45 ps=3.6 w=1.5 l=1
X7 a_2521_2360# Ib.t2 VSS.t4 VSS.t3 sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=1.2 ps=8.6 w=4 l=1
X8 Vout.t2 a_2521_2520.t8 VDD.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.375 pd=2 as=0.375 ps=2 w=1.5 l=1
X9 VDD.t1 a_2521_2520.t9 Vout.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.6 as=0.375 ps=2 w=1.5 l=1
R0 a_2521_2520.n1 a_2521_2520.t4 232.297
R1 a_2521_2520.n0 a_2521_2520.n2 149.061
R2 a_2521_2520.n0 a_2521_2520.t7 97.4272
R3 a_2521_2520.n0 a_2521_2520.t9 96.9802
R4 a_2521_2520.n0 a_2521_2520.t1 96.9791
R5 a_2521_2520.t0 a_2521_2520.n1 91.4315
R6 a_2521_2520.n1 a_2521_2520.t5 96.604
R7 a_2521_2520.n1 a_2521_2520.t3 96.6359
R8 a_2521_2520.n0 a_2521_2520.t8 96.604
R9 a_2521_2520.n2 a_2521_2520.t2 32.8338
R10 a_2521_2520.n2 a_2521_2520.t6 32.8338
R11 a_2521_2520.n1 a_2521_2520.n0 3.00643
R12 VDD.t1 VDD.n16 453.406
R13 VDD.n17 VDD.t1 453.406
R14 VDD.t5 VDD.n29 453.406
R15 VDD.n30 VDD.t5 453.406
R16 VDD.n23 VDD.t4 327.976
R17 VDD.n23 VDD.t0 242.024
R18 VDD.n9 VDD.n8 159.805
R19 VDD.n33 VDD.n32 151.044
R20 VDD.n8 VDD.t2 32.8338
R21 VDD.n8 VDD.t3 32.8338
R22 VDD.n32 VDD.t6 32.8338
R23 VDD.n32 VDD.t7 32.8338
R24 VDD.n15 VDD.n4 27.1064
R25 VDD.n38 VDD.n37 27.1064
R26 VDD.n16 VDD.n5 24.8327
R27 VDD.n18 VDD.n17 24.8327
R28 VDD.n29 VDD.n26 24.8327
R29 VDD.n31 VDD.n30 24.8327
R30 VDD.n34 VDD.n33 12.4943
R31 VDD.n10 VDD.n9 11.8298
R32 VDD.n17 VDD.n4 11.0627
R33 VDD.n16 VDD.n15 11.0627
R34 VDD.n37 VDD.n30 11.0627
R35 VDD.n38 VDD.n29 11.0627
R36 VDD.n37 VDD.n36 9.3005
R37 VDD.n39 VDD.n38 9.3005
R38 VDD.n43 VDD.n42 9.3005
R39 VDD.n41 VDD.n40 9.3005
R40 VDD.n28 VDD.n27 9.3005
R41 VDD.n35 VDD.n34 9.3005
R42 VDD.n10 VDD.n6 9.3005
R43 VDD.n13 VDD.n12 9.3005
R44 VDD.n11 VDD.n3 9.3005
R45 VDD.n7 VDD.n4 9.3005
R46 VDD.n15 VDD.n14 9.3005
R47 VDD.n19 VDD.n2 9.3005
R48 VDD.n21 VDD.n20 9.3005
R49 VDD.n22 VDD.n0 9.3005
R50 VDD.n49 VDD.n48 9.3005
R51 VDD.n47 VDD.n1 9.3005
R52 VDD.n46 VDD.n45 9.3005
R53 VDD.n44 VDD.n25 9.3005
R54 VDD.n24 VDD.n23 8.81002
R55 VDD.n12 VDD.n10 6.58336
R56 VDD.n12 VDD.n11 6.58336
R57 VDD.n11 VDD.n2 6.58336
R58 VDD.n21 VDD.n2 6.58336
R59 VDD.n22 VDD.n21 6.58336
R60 VDD.n48 VDD.n47 6.58336
R61 VDD.n47 VDD.n46 6.58336
R62 VDD.n46 VDD.n25 6.58336
R63 VDD.n42 VDD.n25 6.58336
R64 VDD.n42 VDD.n41 6.58336
R65 VDD.n41 VDD.n27 6.58336
R66 VDD.n34 VDD.n27 6.58336
R67 VDD.n24 VDD.n22 3.29193
R68 VDD.n48 VDD.n24 3.29193
R69 VDD VDD.n50 0.749201
R70 VDD.n20 VDD.n19 0.0647857
R71 VDD.n20 VDD.n0 0.0647857
R72 VDD.n49 VDD.n1 0.0647857
R73 VDD.n45 VDD.n1 0.0647857
R74 VDD.n45 VDD.n44 0.0647857
R75 VDD.n44 VDD.n43 0.0527783
R76 VDD.n50 VDD.n0 0.0326429
R77 VDD.n50 VDD.n49 0.0326429
R78 VDD.n40 VDD.n26 0.0302414
R79 VDD.n39 VDD.n28 0.0302414
R80 VDD.n36 VDD.n35 0.0302414
R81 VDD.n14 VDD.n6 0.0173103
R82 VDD.n13 VDD.n7 0.0173103
R83 VDD.n18 VDD.n3 0.0173103
R84 VDD.n19 VDD.n18 0.0165714
R85 VDD.n6 VDD.n5 0.0147241
R86 VDD.n14 VDD.n13 0.0147241
R87 VDD.n7 VDD.n3 0.0147241
R88 VDD.n33 VDD.n31 0.013
R89 VDD.n9 VDD.n5 0.013
R90 VDD.n43 VDD.n26 0.0017931
R91 VDD.n40 VDD.n39 0.0017931
R92 VDD.n36 VDD.n28 0.0017931
R93 VDD.n35 VDD.n31 0.0017931
R94 Vp Vp.t0 343.64
R95 VSS.n325 VSS.n94 2346.67
R96 VSS.n326 VSS.n325 2346.67
R97 VSS.n327 VSS.n326 2346.67
R98 VSS.n327 VSS.n88 2346.67
R99 VSS.n335 VSS.n88 2346.67
R100 VSS.n336 VSS.n335 2346.67
R101 VSS.n337 VSS.n336 2346.67
R102 VSS.n337 VSS.n82 2346.67
R103 VSS.n345 VSS.n82 2346.67
R104 VSS.n346 VSS.n345 2346.67
R105 VSS.n347 VSS.n346 2346.67
R106 VSS.n347 VSS.n76 2346.67
R107 VSS.n355 VSS.n76 2346.67
R108 VSS.n356 VSS.n355 2346.67
R109 VSS.n357 VSS.n356 2346.67
R110 VSS.n357 VSS.n70 2346.67
R111 VSS.n365 VSS.n70 2346.67
R112 VSS.n366 VSS.n365 2346.67
R113 VSS.n367 VSS.n366 2346.67
R114 VSS.n367 VSS.n64 2346.67
R115 VSS.n375 VSS.n64 2346.67
R116 VSS.n317 VSS.n316 2236.46
R117 VSS.n377 VSS.n376 1994.09
R118 VSS.n316 VSS.n315 1750.28
R119 VSS.n315 VSS.n100 1750.28
R120 VSS.n187 VSS.n100 1750.28
R121 VSS.n188 VSS.n187 1750.28
R122 VSS.n189 VSS.n188 1750.28
R123 VSS.n191 VSS.n189 1750.28
R124 VSS.n192 VSS.n191 1750.28
R125 VSS.n193 VSS.n192 1750.28
R126 VSS.n194 VSS.n193 1750.28
R127 VSS.n196 VSS.n194 1750.28
R128 VSS.n197 VSS.n196 1750.28
R129 VSS.n198 VSS.n197 1750.28
R130 VSS.n199 VSS.n198 1750.28
R131 VSS.n201 VSS.n199 1750.28
R132 VSS.n202 VSS.n201 1750.28
R133 VSS.n203 VSS.n202 1750.28
R134 VSS.n204 VSS.n203 1750.28
R135 VSS.n377 VSS.n58 1560.59
R136 VSS.n385 VSS.n58 1560.59
R137 VSS.n386 VSS.n385 1560.59
R138 VSS.n387 VSS.n386 1560.59
R139 VSS.n387 VSS.n52 1560.59
R140 VSS.n395 VSS.n52 1560.59
R141 VSS.n396 VSS.n395 1560.59
R142 VSS.n397 VSS.n396 1560.59
R143 VSS.n397 VSS.n46 1560.59
R144 VSS.n405 VSS.n46 1560.59
R145 VSS.n406 VSS.n405 1560.59
R146 VSS.n407 VSS.n406 1560.59
R147 VSS.n407 VSS.n40 1560.59
R148 VSS.n415 VSS.n40 1560.59
R149 VSS.n416 VSS.n415 1560.59
R150 VSS.n417 VSS.n416 1560.59
R151 VSS.n417 VSS.n21 1560.59
R152 VSS.n317 VSS.n94 1140.74
R153 VSS.n318 VSS.n317 1046.88
R154 VSS.n376 VSS.n63 996.823
R155 VSS.n318 VSS.n99 783.717
R156 VSS.n378 VSS.n63 783.717
R157 VSS.n494 VSS.n493 783.717
R158 VSS.n182 VSS.n154 783.717
R159 VSS.n99 VSS.n98 585
R160 VSS.n316 VSS.n99 585
R161 VSS.n314 VSS.n313 585
R162 VSS.n315 VSS.n314 585
R163 VSS.n102 VSS.n101 585
R164 VSS.n101 VSS.n100 585
R165 VSS.n309 VSS.n104 585
R166 VSS.n187 VSS.n104 585
R167 VSS.n308 VSS.n105 585
R168 VSS.n188 VSS.n105 585
R169 VSS.n307 VSS.n106 585
R170 VSS.n189 VSS.n106 585
R171 VSS.n190 VSS.n107 585
R172 VSS.n191 VSS.n190 585
R173 VSS.n303 VSS.n109 585
R174 VSS.n192 VSS.n109 585
R175 VSS.n302 VSS.n110 585
R176 VSS.n193 VSS.n110 585
R177 VSS.n301 VSS.n111 585
R178 VSS.n194 VSS.n111 585
R179 VSS.n195 VSS.n112 585
R180 VSS.n196 VSS.n195 585
R181 VSS.n297 VSS.n114 585
R182 VSS.n197 VSS.n114 585
R183 VSS.n296 VSS.n115 585
R184 VSS.n198 VSS.n115 585
R185 VSS.n295 VSS.n116 585
R186 VSS.n199 VSS.n116 585
R187 VSS.n200 VSS.n117 585
R188 VSS.n201 VSS.n200 585
R189 VSS.n291 VSS.n119 585
R190 VSS.n202 VSS.n119 585
R191 VSS.n290 VSS.n120 585
R192 VSS.n203 VSS.n120 585
R193 VSS.n289 VSS.n121 585
R194 VSS.n204 VSS.n121 585
R195 VSS.n184 VSS.n122 585
R196 VSS.n285 VSS.n124 585
R197 VSS.n284 VSS.n125 585
R198 VSS.n186 VSS.n125 585
R199 VSS.n283 VSS.n126 585
R200 VSS.n167 VSS.n127 585
R201 VSS.n279 VSS.n129 585
R202 VSS.n278 VSS.n130 585
R203 VSS.n277 VSS.n131 585
R204 VSS.n170 VSS.n132 585
R205 VSS.n273 VSS.n134 585
R206 VSS.n272 VSS.n135 585
R207 VSS.n271 VSS.n136 585
R208 VSS.n173 VSS.n137 585
R209 VSS.n267 VSS.n139 585
R210 VSS.n266 VSS.n140 585
R211 VSS.n265 VSS.n141 585
R212 VSS.n176 VSS.n142 585
R213 VSS.n261 VSS.n144 585
R214 VSS.n260 VSS.n145 585
R215 VSS.n259 VSS.n146 585
R216 VSS.n179 VSS.n147 585
R217 VSS.n255 VSS.n149 585
R218 VSS.n254 VSS.n150 585
R219 VSS.n253 VSS.n151 585
R220 VSS.n182 VSS.n152 585
R221 VSS.n319 VSS.n318 585
R222 VSS.n96 VSS.n95 585
R223 VSS.n95 VSS.n94 585
R224 VSS.n324 VSS.n323 585
R225 VSS.n325 VSS.n324 585
R226 VSS.n93 VSS.n92 585
R227 VSS.n326 VSS.n93 585
R228 VSS.n329 VSS.n328 585
R229 VSS.n328 VSS.n327 585
R230 VSS.n90 VSS.n89 585
R231 VSS.n89 VSS.n88 585
R232 VSS.n334 VSS.n333 585
R233 VSS.n335 VSS.n334 585
R234 VSS.n87 VSS.n86 585
R235 VSS.n336 VSS.n87 585
R236 VSS.n339 VSS.n338 585
R237 VSS.n338 VSS.n337 585
R238 VSS.n84 VSS.n83 585
R239 VSS.n83 VSS.n82 585
R240 VSS.n344 VSS.n343 585
R241 VSS.n345 VSS.n344 585
R242 VSS.n81 VSS.n80 585
R243 VSS.n346 VSS.n81 585
R244 VSS.n349 VSS.n348 585
R245 VSS.n348 VSS.n347 585
R246 VSS.n78 VSS.n77 585
R247 VSS.n77 VSS.n76 585
R248 VSS.n354 VSS.n353 585
R249 VSS.n355 VSS.n354 585
R250 VSS.n75 VSS.n74 585
R251 VSS.n356 VSS.n75 585
R252 VSS.n359 VSS.n358 585
R253 VSS.n358 VSS.n357 585
R254 VSS.n72 VSS.n71 585
R255 VSS.n71 VSS.n70 585
R256 VSS.n364 VSS.n363 585
R257 VSS.n365 VSS.n364 585
R258 VSS.n69 VSS.n68 585
R259 VSS.n366 VSS.n69 585
R260 VSS.n369 VSS.n368 585
R261 VSS.n368 VSS.n367 585
R262 VSS.n66 VSS.n65 585
R263 VSS.n65 VSS.n64 585
R264 VSS.n374 VSS.n373 585
R265 VSS.n375 VSS.n374 585
R266 VSS.n63 VSS.n62 585
R267 VSS.n495 VSS.n494 585
R268 VSS.n452 VSS.n18 585
R269 VSS.n454 VSS.n453 585
R270 VSS.n451 VSS.n450 585
R271 VSS.n458 VSS.n449 585
R272 VSS.n459 VSS.n448 585
R273 VSS.n460 VSS.n447 585
R274 VSS.n445 VSS.n444 585
R275 VSS.n464 VSS.n443 585
R276 VSS.n465 VSS.n442 585
R277 VSS.n466 VSS.n441 585
R278 VSS.n439 VSS.n438 585
R279 VSS.n470 VSS.n437 585
R280 VSS.n471 VSS.n436 585
R281 VSS.n472 VSS.n435 585
R282 VSS.n433 VSS.n432 585
R283 VSS.n476 VSS.n431 585
R284 VSS.n477 VSS.n430 585
R285 VSS.n478 VSS.n429 585
R286 VSS.n427 VSS.n426 585
R287 VSS.n482 VSS.n425 585
R288 VSS.n483 VSS.n424 585
R289 VSS.n484 VSS.n423 585
R290 VSS.n36 VSS.n34 585
R291 VSS.n489 VSS.n488 585
R292 VSS.n490 VSS.n489 585
R293 VSS.n35 VSS.n33 585
R294 VSS.n33 VSS.n21 585
R295 VSS.n419 VSS.n418 585
R296 VSS.n418 VSS.n417 585
R297 VSS.n39 VSS.n38 585
R298 VSS.n416 VSS.n39 585
R299 VSS.n414 VSS.n413 585
R300 VSS.n415 VSS.n414 585
R301 VSS.n42 VSS.n41 585
R302 VSS.n41 VSS.n40 585
R303 VSS.n409 VSS.n408 585
R304 VSS.n408 VSS.n407 585
R305 VSS.n45 VSS.n44 585
R306 VSS.n406 VSS.n45 585
R307 VSS.n404 VSS.n403 585
R308 VSS.n405 VSS.n404 585
R309 VSS.n48 VSS.n47 585
R310 VSS.n47 VSS.n46 585
R311 VSS.n399 VSS.n398 585
R312 VSS.n398 VSS.n397 585
R313 VSS.n51 VSS.n50 585
R314 VSS.n396 VSS.n51 585
R315 VSS.n394 VSS.n393 585
R316 VSS.n395 VSS.n394 585
R317 VSS.n54 VSS.n53 585
R318 VSS.n53 VSS.n52 585
R319 VSS.n389 VSS.n388 585
R320 VSS.n388 VSS.n387 585
R321 VSS.n57 VSS.n56 585
R322 VSS.n386 VSS.n57 585
R323 VSS.n384 VSS.n383 585
R324 VSS.n385 VSS.n384 585
R325 VSS.n60 VSS.n59 585
R326 VSS.n59 VSS.n58 585
R327 VSS.n379 VSS.n378 585
R328 VSS.n378 VSS.n377 585
R329 VSS.n493 VSS.n16 585
R330 VSS.n493 VSS.n492 585
R331 VSS.n499 VSS.n15 585
R332 VSS.n20 VSS.n15 585
R333 VSS.n500 VSS.n14 585
R334 VSS.n218 VSS.n14 585
R335 VSS.n501 VSS.n13 585
R336 VSS.n219 VSS.n13 585
R337 VSS.n220 VSS.n11 585
R338 VSS.n221 VSS.n220 585
R339 VSS.n505 VSS.n10 585
R340 VSS.n222 VSS.n10 585
R341 VSS.n506 VSS.n9 585
R342 VSS.n223 VSS.n9 585
R343 VSS.n507 VSS.n8 585
R344 VSS.n224 VSS.n8 585
R345 VSS.n225 VSS.n6 585
R346 VSS.n226 VSS.n225 585
R347 VSS.n512 VSS.n5 585
R348 VSS.n227 VSS.n5 585
R349 VSS.n513 VSS.n4 585
R350 VSS.n228 VSS.n4 585
R351 VSS.n514 VSS.n3 585
R352 VSS.n229 VSS.n3 585
R353 VSS.n166 VSS.n2 585
R354 VSS.n230 VSS.n166 585
R355 VSS.n233 VSS.n232 585
R356 VSS.n232 VSS.n231 585
R357 VSS.n236 VSS.n165 585
R358 VSS.n217 VSS.n165 585
R359 VSS.n237 VSS.n164 585
R360 VSS.n216 VSS.n164 585
R361 VSS.n214 VSS.n162 585
R362 VSS.n215 VSS.n214 585
R363 VSS.n241 VSS.n161 585
R364 VSS.n213 VSS.n161 585
R365 VSS.n242 VSS.n160 585
R366 VSS.n212 VSS.n160 585
R367 VSS.n243 VSS.n159 585
R368 VSS.n211 VSS.n159 585
R369 VSS.n209 VSS.n157 585
R370 VSS.n210 VSS.n209 585
R371 VSS.n247 VSS.n156 585
R372 VSS.n208 VSS.n156 585
R373 VSS.n248 VSS.n155 585
R374 VSS.n207 VSS.n155 585
R375 VSS.n249 VSS.n154 585
R376 VSS.n206 VSS.n154 585
R377 VSS.n376 VSS.n375 423.704
R378 VSS.n318 VSS.n95 308.349
R379 VSS.n324 VSS.n95 308.349
R380 VSS.n324 VSS.n93 308.349
R381 VSS.n328 VSS.n93 308.349
R382 VSS.n328 VSS.n89 308.349
R383 VSS.n334 VSS.n89 308.349
R384 VSS.n334 VSS.n87 308.349
R385 VSS.n338 VSS.n87 308.349
R386 VSS.n338 VSS.n83 308.349
R387 VSS.n344 VSS.n83 308.349
R388 VSS.n344 VSS.n81 308.349
R389 VSS.n348 VSS.n81 308.349
R390 VSS.n348 VSS.n77 308.349
R391 VSS.n354 VSS.n77 308.349
R392 VSS.n354 VSS.n75 308.349
R393 VSS.n358 VSS.n75 308.349
R394 VSS.n358 VSS.n71 308.349
R395 VSS.n364 VSS.n71 308.349
R396 VSS.n364 VSS.n69 308.349
R397 VSS.n368 VSS.n69 308.349
R398 VSS.n368 VSS.n65 308.349
R399 VSS.n374 VSS.n65 308.349
R400 VSS.n374 VSS.n63 308.349
R401 VSS.n378 VSS.n59 308.349
R402 VSS.n384 VSS.n59 308.349
R403 VSS.n384 VSS.n57 308.349
R404 VSS.n388 VSS.n57 308.349
R405 VSS.n388 VSS.n53 308.349
R406 VSS.n394 VSS.n53 308.349
R407 VSS.n394 VSS.n51 308.349
R408 VSS.n398 VSS.n51 308.349
R409 VSS.n398 VSS.n47 308.349
R410 VSS.n404 VSS.n47 308.349
R411 VSS.n404 VSS.n45 308.349
R412 VSS.n408 VSS.n45 308.349
R413 VSS.n408 VSS.n41 308.349
R414 VSS.n414 VSS.n41 308.349
R415 VSS.n414 VSS.n39 308.349
R416 VSS.n418 VSS.n39 308.349
R417 VSS.n418 VSS.n33 308.349
R418 VSS.n489 VSS.n33 308.349
R419 VSS.n489 VSS.n34 308.349
R420 VSS.n424 VSS.n423 308.349
R421 VSS.n426 VSS.n425 308.349
R422 VSS.n430 VSS.n429 308.349
R423 VSS.n432 VSS.n431 308.349
R424 VSS.n436 VSS.n435 308.349
R425 VSS.n438 VSS.n437 308.349
R426 VSS.n442 VSS.n441 308.349
R427 VSS.n444 VSS.n443 308.349
R428 VSS.n448 VSS.n447 308.349
R429 VSS.n450 VSS.n449 308.349
R430 VSS.n453 VSS.n452 308.349
R431 VSS.n155 VSS.n154 308.349
R432 VSS.n156 VSS.n155 308.349
R433 VSS.n209 VSS.n156 308.349
R434 VSS.n209 VSS.n159 308.349
R435 VSS.n160 VSS.n159 308.349
R436 VSS.n161 VSS.n160 308.349
R437 VSS.n214 VSS.n161 308.349
R438 VSS.n214 VSS.n164 308.349
R439 VSS.n165 VSS.n164 308.349
R440 VSS.n232 VSS.n165 308.349
R441 VSS.n232 VSS.n166 308.349
R442 VSS.n166 VSS.n3 308.349
R443 VSS.n4 VSS.n3 308.349
R444 VSS.n5 VSS.n4 308.349
R445 VSS.n225 VSS.n5 308.349
R446 VSS.n225 VSS.n8 308.349
R447 VSS.n9 VSS.n8 308.349
R448 VSS.n10 VSS.n9 308.349
R449 VSS.n220 VSS.n10 308.349
R450 VSS.n220 VSS.n13 308.349
R451 VSS.n14 VSS.n13 308.349
R452 VSS.n15 VSS.n14 308.349
R453 VSS.n493 VSS.n15 308.349
R454 VSS.n314 VSS.n99 308.349
R455 VSS.n314 VSS.n101 308.349
R456 VSS.n104 VSS.n101 308.349
R457 VSS.n105 VSS.n104 308.349
R458 VSS.n106 VSS.n105 308.349
R459 VSS.n190 VSS.n106 308.349
R460 VSS.n190 VSS.n109 308.349
R461 VSS.n110 VSS.n109 308.349
R462 VSS.n111 VSS.n110 308.349
R463 VSS.n195 VSS.n111 308.349
R464 VSS.n195 VSS.n114 308.349
R465 VSS.n115 VSS.n114 308.349
R466 VSS.n116 VSS.n115 308.349
R467 VSS.n200 VSS.n116 308.349
R468 VSS.n200 VSS.n119 308.349
R469 VSS.n120 VSS.n119 308.349
R470 VSS.n121 VSS.n120 308.349
R471 VSS.n184 VSS.n121 308.349
R472 VSS.n125 VSS.n124 308.349
R473 VSS.n126 VSS.n125 308.349
R474 VSS.n167 VSS.n129 308.349
R475 VSS.n131 VSS.n130 308.349
R476 VSS.n170 VSS.n134 308.349
R477 VSS.n136 VSS.n135 308.349
R478 VSS.n173 VSS.n139 308.349
R479 VSS.n141 VSS.n140 308.349
R480 VSS.n176 VSS.n144 308.349
R481 VSS.n146 VSS.n145 308.349
R482 VSS.n179 VSS.n149 308.349
R483 VSS.n151 VSS.n150 308.349
R484 VSS.n205 VSS.n204 267.404
R485 VSS.n491 VSS.n21 238.424
R486 VSS.n186 VSS.n185 231.493
R487 VSS.n186 VSS.n168 231.493
R488 VSS.n186 VSS.n169 231.493
R489 VSS.n186 VSS.n171 231.493
R490 VSS.n186 VSS.n172 231.493
R491 VSS.n186 VSS.n174 231.493
R492 VSS.n186 VSS.n175 231.493
R493 VSS.n186 VSS.n177 231.493
R494 VSS.n186 VSS.n178 231.493
R495 VSS.n186 VSS.n180 231.493
R496 VSS.n186 VSS.n181 231.493
R497 VSS.n186 VSS.n183 231.493
R498 VSS.n490 VSS.n19 231.493
R499 VSS.n490 VSS.n22 231.493
R500 VSS.n490 VSS.n23 231.493
R501 VSS.n490 VSS.n24 231.493
R502 VSS.n490 VSS.n25 231.493
R503 VSS.n490 VSS.n26 231.493
R504 VSS.n490 VSS.n27 231.493
R505 VSS.n490 VSS.n28 231.493
R506 VSS.n490 VSS.n29 231.493
R507 VSS.n490 VSS.n30 231.493
R508 VSS.n490 VSS.n31 231.493
R509 VSS.n490 VSS.n32 231.493
R510 VSS.n207 VSS.n206 162.546
R511 VSS.n208 VSS.n207 162.546
R512 VSS.n210 VSS.n208 162.546
R513 VSS.n211 VSS.n210 162.546
R514 VSS.n212 VSS.n211 162.546
R515 VSS.n215 VSS.n213 162.546
R516 VSS.n216 VSS.n215 162.546
R517 VSS.n217 VSS.n216 162.546
R518 VSS.n231 VSS.n217 162.546
R519 VSS.n231 VSS.n230 162.546
R520 VSS.n230 VSS.n229 162.546
R521 VSS.n229 VSS.n228 162.546
R522 VSS.n228 VSS.n227 162.546
R523 VSS.n227 VSS.n226 162.546
R524 VSS.n226 VSS.n224 162.546
R525 VSS.n222 VSS.n221 162.546
R526 VSS.n221 VSS.n219 162.546
R527 VSS.n219 VSS.n218 162.546
R528 VSS.n218 VSS.n20 162.546
R529 VSS.n492 VSS.n20 162.546
R530 VSS.n224 VSS.t0 155.773
R531 VSS.t2 VSS.n212 142.227
R532 VSS.n423 VSS.n32 122.017
R533 VSS.n425 VSS.n31 122.017
R534 VSS.n429 VSS.n30 122.017
R535 VSS.n431 VSS.n29 122.017
R536 VSS.n435 VSS.n28 122.017
R537 VSS.n437 VSS.n27 122.017
R538 VSS.n441 VSS.n26 122.017
R539 VSS.n443 VSS.n25 122.017
R540 VSS.n447 VSS.n24 122.017
R541 VSS.n449 VSS.n23 122.017
R542 VSS.n453 VSS.n22 122.017
R543 VSS.n494 VSS.n19 122.017
R544 VSS.n185 VSS.n184 122.017
R545 VSS.n168 VSS.n126 122.017
R546 VSS.n169 VSS.n129 122.017
R547 VSS.n171 VSS.n131 122.017
R548 VSS.n172 VSS.n134 122.017
R549 VSS.n174 VSS.n136 122.017
R550 VSS.n175 VSS.n139 122.017
R551 VSS.n177 VSS.n141 122.017
R552 VSS.n178 VSS.n144 122.017
R553 VSS.n180 VSS.n146 122.017
R554 VSS.n181 VSS.n149 122.017
R555 VSS.n183 VSS.n151 122.017
R556 VSS.n185 VSS.n124 122.017
R557 VSS.n168 VSS.n167 122.017
R558 VSS.n169 VSS.n130 122.017
R559 VSS.n171 VSS.n170 122.017
R560 VSS.n172 VSS.n135 122.017
R561 VSS.n174 VSS.n173 122.017
R562 VSS.n175 VSS.n140 122.017
R563 VSS.n177 VSS.n176 122.017
R564 VSS.n178 VSS.n145 122.017
R565 VSS.n180 VSS.n179 122.017
R566 VSS.n181 VSS.n150 122.017
R567 VSS.n183 VSS.n182 122.017
R568 VSS.n452 VSS.n19 122.017
R569 VSS.n450 VSS.n22 122.017
R570 VSS.n448 VSS.n23 122.017
R571 VSS.n444 VSS.n24 122.017
R572 VSS.n442 VSS.n25 122.017
R573 VSS.n438 VSS.n26 122.017
R574 VSS.n436 VSS.n27 122.017
R575 VSS.n432 VSS.n28 122.017
R576 VSS.n430 VSS.n29 122.017
R577 VSS.n426 VSS.n30 122.017
R578 VSS.n424 VSS.n31 122.017
R579 VSS.n34 VSS.n32 122.017
R580 VSS.n206 VSS.n205 119.651
R581 VSS.n491 VSS.n490 117.394
R582 VSS.t5 VSS.n222 112.879
R583 VSS.n492 VSS.n491 97.0759
R584 VSS.n205 VSS.n186 94.8183
R585 VSS.n319 VSS.n98 50.9222
R586 VSS.n249 VSS.n152 50.9222
R587 VSS.n379 VSS.n62 50.9222
R588 VSS.n495 VSS.n16 50.9222
R589 VSS.n223 VSS.t5 49.667
R590 VSS.n163 VSS.t4 22.6843
R591 VSS.n510 VSS.t1 22.6843
R592 VSS.n313 VSS.n98 20.0353
R593 VSS.n313 VSS.n102 20.0353
R594 VSS.n309 VSS.n102 20.0353
R595 VSS.n309 VSS.n308 20.0353
R596 VSS.n308 VSS.n307 20.0353
R597 VSS.n307 VSS.n107 20.0353
R598 VSS.n303 VSS.n107 20.0353
R599 VSS.n303 VSS.n302 20.0353
R600 VSS.n302 VSS.n301 20.0353
R601 VSS.n301 VSS.n112 20.0353
R602 VSS.n297 VSS.n112 20.0353
R603 VSS.n297 VSS.n296 20.0353
R604 VSS.n296 VSS.n295 20.0353
R605 VSS.n295 VSS.n117 20.0353
R606 VSS.n291 VSS.n117 20.0353
R607 VSS.n291 VSS.n290 20.0353
R608 VSS.n290 VSS.n289 20.0353
R609 VSS.n289 VSS.n122 20.0353
R610 VSS.n285 VSS.n122 20.0353
R611 VSS.n285 VSS.n284 20.0353
R612 VSS.n284 VSS.n283 20.0353
R613 VSS.n283 VSS.n127 20.0353
R614 VSS.n279 VSS.n127 20.0353
R615 VSS.n279 VSS.n278 20.0353
R616 VSS.n278 VSS.n277 20.0353
R617 VSS.n277 VSS.n132 20.0353
R618 VSS.n273 VSS.n132 20.0353
R619 VSS.n273 VSS.n272 20.0353
R620 VSS.n272 VSS.n271 20.0353
R621 VSS.n271 VSS.n137 20.0353
R622 VSS.n267 VSS.n137 20.0353
R623 VSS.n267 VSS.n266 20.0353
R624 VSS.n266 VSS.n265 20.0353
R625 VSS.n265 VSS.n142 20.0353
R626 VSS.n261 VSS.n142 20.0353
R627 VSS.n261 VSS.n260 20.0353
R628 VSS.n260 VSS.n259 20.0353
R629 VSS.n259 VSS.n147 20.0353
R630 VSS.n255 VSS.n147 20.0353
R631 VSS.n255 VSS.n254 20.0353
R632 VSS.n254 VSS.n253 20.0353
R633 VSS.n253 VSS.n152 20.0353
R634 VSS.n319 VSS.n96 20.0353
R635 VSS.n323 VSS.n96 20.0353
R636 VSS.n323 VSS.n92 20.0353
R637 VSS.n329 VSS.n92 20.0353
R638 VSS.n329 VSS.n90 20.0353
R639 VSS.n333 VSS.n90 20.0353
R640 VSS.n333 VSS.n86 20.0353
R641 VSS.n339 VSS.n86 20.0353
R642 VSS.n339 VSS.n84 20.0353
R643 VSS.n343 VSS.n84 20.0353
R644 VSS.n343 VSS.n80 20.0353
R645 VSS.n349 VSS.n80 20.0353
R646 VSS.n349 VSS.n78 20.0353
R647 VSS.n353 VSS.n78 20.0353
R648 VSS.n353 VSS.n74 20.0353
R649 VSS.n359 VSS.n74 20.0353
R650 VSS.n359 VSS.n72 20.0353
R651 VSS.n363 VSS.n72 20.0353
R652 VSS.n363 VSS.n68 20.0353
R653 VSS.n369 VSS.n68 20.0353
R654 VSS.n369 VSS.n66 20.0353
R655 VSS.n373 VSS.n66 20.0353
R656 VSS.n373 VSS.n62 20.0353
R657 VSS.n379 VSS.n60 20.0353
R658 VSS.n383 VSS.n60 20.0353
R659 VSS.n383 VSS.n56 20.0353
R660 VSS.n389 VSS.n56 20.0353
R661 VSS.n389 VSS.n54 20.0353
R662 VSS.n393 VSS.n54 20.0353
R663 VSS.n393 VSS.n50 20.0353
R664 VSS.n399 VSS.n50 20.0353
R665 VSS.n399 VSS.n48 20.0353
R666 VSS.n403 VSS.n48 20.0353
R667 VSS.n403 VSS.n44 20.0353
R668 VSS.n409 VSS.n44 20.0353
R669 VSS.n409 VSS.n42 20.0353
R670 VSS.n413 VSS.n42 20.0353
R671 VSS.n413 VSS.n38 20.0353
R672 VSS.n419 VSS.n38 20.0353
R673 VSS.n419 VSS.n35 20.0353
R674 VSS.n488 VSS.n35 20.0353
R675 VSS.n488 VSS.n36 20.0353
R676 VSS.n484 VSS.n36 20.0353
R677 VSS.n484 VSS.n483 20.0353
R678 VSS.n483 VSS.n482 20.0353
R679 VSS.n482 VSS.n427 20.0353
R680 VSS.n478 VSS.n427 20.0353
R681 VSS.n478 VSS.n477 20.0353
R682 VSS.n477 VSS.n476 20.0353
R683 VSS.n476 VSS.n433 20.0353
R684 VSS.n472 VSS.n433 20.0353
R685 VSS.n472 VSS.n471 20.0353
R686 VSS.n471 VSS.n470 20.0353
R687 VSS.n470 VSS.n439 20.0353
R688 VSS.n466 VSS.n439 20.0353
R689 VSS.n466 VSS.n465 20.0353
R690 VSS.n465 VSS.n464 20.0353
R691 VSS.n464 VSS.n445 20.0353
R692 VSS.n460 VSS.n445 20.0353
R693 VSS.n460 VSS.n459 20.0353
R694 VSS.n459 VSS.n458 20.0353
R695 VSS.n458 VSS.n451 20.0353
R696 VSS.n454 VSS.n451 20.0353
R697 VSS.n454 VSS.n18 20.0353
R698 VSS.n495 VSS.n18 20.0353
R699 VSS.n249 VSS.n248 20.0353
R700 VSS.n248 VSS.n247 20.0353
R701 VSS.n247 VSS.n157 20.0353
R702 VSS.n243 VSS.n157 20.0353
R703 VSS.n243 VSS.n242 20.0353
R704 VSS.n242 VSS.n241 20.0353
R705 VSS.n241 VSS.n162 20.0353
R706 VSS.n237 VSS.n162 20.0353
R707 VSS.n237 VSS.n236 20.0353
R708 VSS.n236 VSS.n233 20.0353
R709 VSS.n233 VSS.n2 20.0353
R710 VSS.n514 VSS.n2 20.0353
R711 VSS.n514 VSS.n513 20.0353
R712 VSS.n513 VSS.n512 20.0353
R713 VSS.n512 VSS.n6 20.0353
R714 VSS.n507 VSS.n6 20.0353
R715 VSS.n507 VSS.n506 20.0353
R716 VSS.n506 VSS.n505 20.0353
R717 VSS.n505 VSS.n11 20.0353
R718 VSS.n501 VSS.n11 20.0353
R719 VSS.n501 VSS.n500 20.0353
R720 VSS.n500 VSS.n499 20.0353
R721 VSS.n499 VSS.n16 20.0353
R722 VSS.t3 VSS.t2 13.5459
R723 VSS.n497 VSS.n16 9.3005
R724 VSS.n499 VSS.n498 9.3005
R725 VSS.n496 VSS.n495 9.3005
R726 VSS.n18 VSS.n17 9.3005
R727 VSS.n455 VSS.n454 9.3005
R728 VSS.n456 VSS.n451 9.3005
R729 VSS.n458 VSS.n457 9.3005
R730 VSS.n459 VSS.n446 9.3005
R731 VSS.n461 VSS.n460 9.3005
R732 VSS.n462 VSS.n445 9.3005
R733 VSS.n464 VSS.n463 9.3005
R734 VSS.n465 VSS.n440 9.3005
R735 VSS.n467 VSS.n466 9.3005
R736 VSS.n468 VSS.n439 9.3005
R737 VSS.n470 VSS.n469 9.3005
R738 VSS.n471 VSS.n434 9.3005
R739 VSS.n473 VSS.n472 9.3005
R740 VSS.n474 VSS.n433 9.3005
R741 VSS.n476 VSS.n475 9.3005
R742 VSS.n477 VSS.n428 9.3005
R743 VSS.n479 VSS.n478 9.3005
R744 VSS.n480 VSS.n427 9.3005
R745 VSS.n482 VSS.n481 9.3005
R746 VSS.n483 VSS.n422 9.3005
R747 VSS.n485 VSS.n484 9.3005
R748 VSS.n486 VSS.n36 9.3005
R749 VSS.n488 VSS.n487 9.3005
R750 VSS.n421 VSS.n35 9.3005
R751 VSS.n420 VSS.n419 9.3005
R752 VSS.n38 VSS.n37 9.3005
R753 VSS.n413 VSS.n412 9.3005
R754 VSS.n411 VSS.n42 9.3005
R755 VSS.n410 VSS.n409 9.3005
R756 VSS.n44 VSS.n43 9.3005
R757 VSS.n403 VSS.n402 9.3005
R758 VSS.n401 VSS.n48 9.3005
R759 VSS.n400 VSS.n399 9.3005
R760 VSS.n50 VSS.n49 9.3005
R761 VSS.n393 VSS.n392 9.3005
R762 VSS.n391 VSS.n54 9.3005
R763 VSS.n390 VSS.n389 9.3005
R764 VSS.n56 VSS.n55 9.3005
R765 VSS.n383 VSS.n382 9.3005
R766 VSS.n381 VSS.n60 9.3005
R767 VSS.n380 VSS.n379 9.3005
R768 VSS.n320 VSS.n319 9.3005
R769 VSS.n321 VSS.n96 9.3005
R770 VSS.n323 VSS.n322 9.3005
R771 VSS.n92 VSS.n91 9.3005
R772 VSS.n330 VSS.n329 9.3005
R773 VSS.n331 VSS.n90 9.3005
R774 VSS.n333 VSS.n332 9.3005
R775 VSS.n86 VSS.n85 9.3005
R776 VSS.n340 VSS.n339 9.3005
R777 VSS.n341 VSS.n84 9.3005
R778 VSS.n343 VSS.n342 9.3005
R779 VSS.n80 VSS.n79 9.3005
R780 VSS.n350 VSS.n349 9.3005
R781 VSS.n351 VSS.n78 9.3005
R782 VSS.n353 VSS.n352 9.3005
R783 VSS.n74 VSS.n73 9.3005
R784 VSS.n360 VSS.n359 9.3005
R785 VSS.n361 VSS.n72 9.3005
R786 VSS.n363 VSS.n362 9.3005
R787 VSS.n68 VSS.n67 9.3005
R788 VSS.n370 VSS.n369 9.3005
R789 VSS.n371 VSS.n66 9.3005
R790 VSS.n373 VSS.n372 9.3005
R791 VSS.n62 VSS.n61 9.3005
R792 VSS.n98 VSS.n97 9.3005
R793 VSS.n313 VSS.n312 9.3005
R794 VSS.n311 VSS.n102 9.3005
R795 VSS.n310 VSS.n309 9.3005
R796 VSS.n308 VSS.n103 9.3005
R797 VSS.n307 VSS.n306 9.3005
R798 VSS.n305 VSS.n107 9.3005
R799 VSS.n304 VSS.n303 9.3005
R800 VSS.n302 VSS.n108 9.3005
R801 VSS.n301 VSS.n300 9.3005
R802 VSS.n299 VSS.n112 9.3005
R803 VSS.n298 VSS.n297 9.3005
R804 VSS.n296 VSS.n113 9.3005
R805 VSS.n295 VSS.n294 9.3005
R806 VSS.n293 VSS.n117 9.3005
R807 VSS.n292 VSS.n291 9.3005
R808 VSS.n290 VSS.n118 9.3005
R809 VSS.n289 VSS.n288 9.3005
R810 VSS.n287 VSS.n122 9.3005
R811 VSS.n286 VSS.n285 9.3005
R812 VSS.n284 VSS.n123 9.3005
R813 VSS.n283 VSS.n282 9.3005
R814 VSS.n281 VSS.n127 9.3005
R815 VSS.n280 VSS.n279 9.3005
R816 VSS.n278 VSS.n128 9.3005
R817 VSS.n277 VSS.n276 9.3005
R818 VSS.n275 VSS.n132 9.3005
R819 VSS.n274 VSS.n273 9.3005
R820 VSS.n272 VSS.n133 9.3005
R821 VSS.n271 VSS.n270 9.3005
R822 VSS.n269 VSS.n137 9.3005
R823 VSS.n268 VSS.n267 9.3005
R824 VSS.n266 VSS.n138 9.3005
R825 VSS.n265 VSS.n264 9.3005
R826 VSS.n263 VSS.n142 9.3005
R827 VSS.n262 VSS.n261 9.3005
R828 VSS.n260 VSS.n143 9.3005
R829 VSS.n259 VSS.n258 9.3005
R830 VSS.n257 VSS.n147 9.3005
R831 VSS.n256 VSS.n255 9.3005
R832 VSS.n254 VSS.n148 9.3005
R833 VSS.n253 VSS.n252 9.3005
R834 VSS.n251 VSS.n152 9.3005
R835 VSS.n248 VSS.n153 9.3005
R836 VSS.n250 VSS.n249 9.3005
R837 VSS.n500 VSS.n12 9.3005
R838 VSS.n502 VSS.n501 9.3005
R839 VSS.n503 VSS.n11 9.3005
R840 VSS.n505 VSS.n504 9.3005
R841 VSS.n506 VSS.n7 9.3005
R842 VSS.n508 VSS.n507 9.3005
R843 VSS.n509 VSS.n6 9.3005
R844 VSS.n512 VSS.n511 9.3005
R845 VSS.n513 VSS.n1 9.3005
R846 VSS.n515 VSS.n514 9.3005
R847 VSS.n2 VSS.n0 9.3005
R848 VSS.n234 VSS.n233 9.3005
R849 VSS.n236 VSS.n235 9.3005
R850 VSS.n238 VSS.n237 9.3005
R851 VSS.n239 VSS.n162 9.3005
R852 VSS.n241 VSS.n240 9.3005
R853 VSS.n242 VSS.n158 9.3005
R854 VSS.n244 VSS.n243 9.3005
R855 VSS.n245 VSS.n157 9.3005
R856 VSS.n247 VSS.n246 9.3005
R857 VSS.n213 VSS.t3 6.7732
R858 VSS.t0 VSS.n223 6.7732
R859 VSS VSS.n516 0.747416
R860 VSS.n497 VSS.n496 0.497783
R861 VSS.n380 VSS.n61 0.497783
R862 VSS.n320 VSS.n97 0.497783
R863 VSS.n251 VSS.n250 0.497783
R864 VSS.n498 VSS.n497 0.196152
R865 VSS.n381 VSS.n380 0.196152
R866 VSS.n382 VSS.n381 0.196152
R867 VSS.n382 VSS.n55 0.196152
R868 VSS.n390 VSS.n55 0.196152
R869 VSS.n391 VSS.n390 0.196152
R870 VSS.n392 VSS.n391 0.196152
R871 VSS.n392 VSS.n49 0.196152
R872 VSS.n400 VSS.n49 0.196152
R873 VSS.n401 VSS.n400 0.196152
R874 VSS.n402 VSS.n401 0.196152
R875 VSS.n402 VSS.n43 0.196152
R876 VSS.n410 VSS.n43 0.196152
R877 VSS.n411 VSS.n410 0.196152
R878 VSS.n412 VSS.n411 0.196152
R879 VSS.n412 VSS.n37 0.196152
R880 VSS.n420 VSS.n37 0.196152
R881 VSS.n421 VSS.n420 0.196152
R882 VSS.n487 VSS.n421 0.196152
R883 VSS.n487 VSS.n486 0.196152
R884 VSS.n486 VSS.n485 0.196152
R885 VSS.n485 VSS.n422 0.196152
R886 VSS.n481 VSS.n422 0.196152
R887 VSS.n481 VSS.n480 0.196152
R888 VSS.n480 VSS.n479 0.196152
R889 VSS.n479 VSS.n428 0.196152
R890 VSS.n475 VSS.n428 0.196152
R891 VSS.n475 VSS.n474 0.196152
R892 VSS.n474 VSS.n473 0.196152
R893 VSS.n473 VSS.n434 0.196152
R894 VSS.n469 VSS.n434 0.196152
R895 VSS.n469 VSS.n468 0.196152
R896 VSS.n468 VSS.n467 0.196152
R897 VSS.n467 VSS.n440 0.196152
R898 VSS.n463 VSS.n440 0.196152
R899 VSS.n463 VSS.n462 0.196152
R900 VSS.n462 VSS.n461 0.196152
R901 VSS.n461 VSS.n446 0.196152
R902 VSS.n457 VSS.n446 0.196152
R903 VSS.n457 VSS.n456 0.196152
R904 VSS.n456 VSS.n455 0.196152
R905 VSS.n455 VSS.n17 0.196152
R906 VSS.n496 VSS.n17 0.196152
R907 VSS.n321 VSS.n320 0.196152
R908 VSS.n322 VSS.n321 0.196152
R909 VSS.n322 VSS.n91 0.196152
R910 VSS.n330 VSS.n91 0.196152
R911 VSS.n331 VSS.n330 0.196152
R912 VSS.n332 VSS.n331 0.196152
R913 VSS.n332 VSS.n85 0.196152
R914 VSS.n340 VSS.n85 0.196152
R915 VSS.n341 VSS.n340 0.196152
R916 VSS.n342 VSS.n341 0.196152
R917 VSS.n342 VSS.n79 0.196152
R918 VSS.n350 VSS.n79 0.196152
R919 VSS.n351 VSS.n350 0.196152
R920 VSS.n352 VSS.n351 0.196152
R921 VSS.n352 VSS.n73 0.196152
R922 VSS.n360 VSS.n73 0.196152
R923 VSS.n361 VSS.n360 0.196152
R924 VSS.n362 VSS.n361 0.196152
R925 VSS.n362 VSS.n67 0.196152
R926 VSS.n370 VSS.n67 0.196152
R927 VSS.n371 VSS.n370 0.196152
R928 VSS.n372 VSS.n371 0.196152
R929 VSS.n372 VSS.n61 0.196152
R930 VSS.n312 VSS.n97 0.196152
R931 VSS.n312 VSS.n311 0.196152
R932 VSS.n311 VSS.n310 0.196152
R933 VSS.n310 VSS.n103 0.196152
R934 VSS.n306 VSS.n103 0.196152
R935 VSS.n306 VSS.n305 0.196152
R936 VSS.n305 VSS.n304 0.196152
R937 VSS.n304 VSS.n108 0.196152
R938 VSS.n300 VSS.n108 0.196152
R939 VSS.n300 VSS.n299 0.196152
R940 VSS.n299 VSS.n298 0.196152
R941 VSS.n298 VSS.n113 0.196152
R942 VSS.n294 VSS.n113 0.196152
R943 VSS.n294 VSS.n293 0.196152
R944 VSS.n293 VSS.n292 0.196152
R945 VSS.n292 VSS.n118 0.196152
R946 VSS.n288 VSS.n118 0.196152
R947 VSS.n288 VSS.n287 0.196152
R948 VSS.n287 VSS.n286 0.196152
R949 VSS.n286 VSS.n123 0.196152
R950 VSS.n282 VSS.n123 0.196152
R951 VSS.n282 VSS.n281 0.196152
R952 VSS.n281 VSS.n280 0.196152
R953 VSS.n280 VSS.n128 0.196152
R954 VSS.n276 VSS.n128 0.196152
R955 VSS.n276 VSS.n275 0.196152
R956 VSS.n275 VSS.n274 0.196152
R957 VSS.n274 VSS.n133 0.196152
R958 VSS.n270 VSS.n133 0.196152
R959 VSS.n270 VSS.n269 0.196152
R960 VSS.n269 VSS.n268 0.196152
R961 VSS.n268 VSS.n138 0.196152
R962 VSS.n264 VSS.n138 0.196152
R963 VSS.n264 VSS.n263 0.196152
R964 VSS.n263 VSS.n262 0.196152
R965 VSS.n262 VSS.n143 0.196152
R966 VSS.n258 VSS.n143 0.196152
R967 VSS.n258 VSS.n257 0.196152
R968 VSS.n257 VSS.n256 0.196152
R969 VSS.n256 VSS.n148 0.196152
R970 VSS.n252 VSS.n148 0.196152
R971 VSS.n252 VSS.n251 0.196152
R972 VSS.n250 VSS.n153 0.196152
R973 VSS.n498 VSS.n12 0.108643
R974 VSS.n246 VSS.n153 0.0648884
R975 VSS.n246 VSS.n245 0.0386356
R976 VSS.n245 VSS.n244 0.0386356
R977 VSS.n244 VSS.n158 0.0386356
R978 VSS.n240 VSS.n158 0.0386356
R979 VSS.n240 VSS.n239 0.0386356
R980 VSS.n239 VSS.n238 0.0386356
R981 VSS.n235 VSS.n234 0.0386356
R982 VSS.n234 VSS.n0 0.0386356
R983 VSS.n515 VSS.n1 0.0386356
R984 VSS.n511 VSS.n1 0.0386356
R985 VSS.n509 VSS.n508 0.0386356
R986 VSS.n508 VSS.n7 0.0386356
R987 VSS.n504 VSS.n7 0.0386356
R988 VSS.n504 VSS.n503 0.0386356
R989 VSS.n503 VSS.n502 0.0386356
R990 VSS.n502 VSS.n12 0.0386356
R991 VSS.n235 VSS.n163 0.0354576
R992 VSS.n511 VSS.n510 0.0322797
R993 VSS.n516 VSS.n515 0.0248644
R994 VSS.n516 VSS.n0 0.0142712
R995 VSS.n510 VSS.n509 0.00685593
R996 VSS.n238 VSS.n163 0.00367797
R997 Vn Vn.t0 342.793
R998 Vout.n1 Vout.t3 232.304
R999 Vout.n1 Vout.n0 151.816
R1000 Vout.n2 Vout.t0 91.2896
R1001 Vout.n0 Vout.t1 32.8338
R1002 Vout.n0 Vout.t2 32.8338
R1003 Vout Vout.n2 1.18443
R1004 Vout.n2 Vout.n1 0.140437
R1005 Ib.n4 Ib.n3 184.74
R1006 Ib.n7 Ib.t2 157.993
R1007 Ib.n4 Ib.t0 96.4005
R1008 Ib.n5 Ib.n4 77.1778
R1009 Ib.n3 Ib.n1 27.1064
R1010 Ib.n6 Ib.n5 23.0638
R1011 Ib.n2 Ib.t1 22.9674
R1012 Ib.n5 Ib.n1 11.3247
R1013 Ib.n1 Ib.n0 9.3005
R1014 Ib.n3 Ib.n2 9.3005
R1015 Ib Ib.n7 1.87558
R1016 Ib.n7 Ib.n6 0.848326
R1017 Ib.n6 Ib.n0 0.196152
R1018 Ib.n2 Ib.n0 0.196152
C0 a_2521_2360# Vout 0.257311f
C1 Vp VDD 0.017362f
C2 a_2521_2360# VDD 0.015449f
C3 Ib Vp 0.089627f
C4 Ib a_2521_2360# 0.480542f
C5 VDD Vout 0.672888f
C6 Vp Vn 0.024179f
C7 Vn a_2521_2360# 0.129522f
C8 Vp a_2521_2360# 0.214004f
C9 Vn Vout 0.08263f
C10 Vn VDD 0.023571f
C11 Ib VSS 2.51866f
C12 Vn VSS 0.53857f
C13 Vp VSS 0.576004f
C14 Vout VSS 0.503831f
C15 VDD VSS 7.53227f
C16 a_2521_2360# VSS 1.13762f
C17 VDD.n5 VSS 0.010806f
C18 VDD.n8 VSS 0.017963f
C19 VDD.n9 VSS 0.149115f
C20 VDD.n10 VSS 0.017578f
C21 VDD.t1 VSS 0.01136f
C22 VDD.n18 VSS 0.012592f
C23 VDD.t0 VSS 0.746478f
C24 VDD.t4 VSS 0.677795f
C25 VDD.n23 VSS 0.357206f
C26 VDD.n24 VSS -0.093452f
C27 VDD.n26 VSS 0.012193f
C28 VDD.t5 VSS 0.01136f
C29 VDD.n32 VSS 0.015111f
C30 VDD.n33 VSS 0.097393f
C31 VDD.n34 VSS 0.017489f
C32 VDD.n50 VSS 0.131514f
C33 a_2521_2520.n0 VSS 0.597736f
C34 a_2521_2520.n1 VSS 0.661915f
C35 a_2521_2520.t3 VSS 0.193837f
C36 a_2521_2520.t5 VSS 0.19382f
C37 a_2521_2520.t1 VSS 0.194155f
C38 a_2521_2520.t9 VSS 0.194156f
C39 a_2521_2520.t8 VSS 0.19382f
C40 a_2521_2520.t7 VSS 0.194751f
C41 a_2521_2520.t2 VSS 0.02487f
C42 a_2521_2520.t6 VSS 0.02487f
C43 a_2521_2520.n2 VSS 0.050484f
C44 a_2521_2520.t4 VSS 0.040067f
C45 a_2521_2520.t0 VSS 0.035518f
.ends

